module ctrl (
    input [2:0] funct3,
    input [6:0] funct7,
    input [6:0] opcode,
    input zero,
    output pc_src,
    output result_src,
    output mem_write,
    output [1:0] alu_op,
    output alu_src,
    output [1:0] imm_src,
    output reg_write
);


    
endmodule